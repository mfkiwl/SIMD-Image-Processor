library verilog;
use verilog.vl_types.all;
entity tb_lab6 is
end tb_lab6;
